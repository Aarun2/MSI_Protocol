module cache_core();

    input clk, rst_n, rd;
    input [:0] wr_data;
    input [:0] wr_addr, rd_addr;
    output rd_data;
    output rd_rdy, wr_rdy;



endmodule